library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package gen_pkg is
	subtype myvec is std_logic_vector(1 downto 0);
end package gen_pkg;
